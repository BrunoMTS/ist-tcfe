T1_CIRCUIT

R1 n1 n2 1.03034608494k
R2 n2 n3 2.03076273175k
R3 n2 n5 3.09442618781k
R4 GND n5 4.08713017488k
R5 n4 n5 3.00518812223k
R6 n6a n6 2.03106965039k
R7 n6 n7 1.04759435052k
VO GND n6a dc 0
Va n1 GND dc 5.01015797903
Id n7 n4 dc 1.02637626609m
Hc n5 n7 VO 8.13697715515k
Gb n4 n3 n2 n5 7.27607852163m
.op
.end

